
module hex7
(
    input  wire [3:0] i, // Вход
    output wire [6:0] o  // Выход
);

assign o = (
    //                6543210
    i == 4'b0000 ? 7'b1000000 : // 0
    i == 4'b0001 ? 7'b1111001 : // 1
    i == 4'b0010 ? 7'b0100100 : // 2
    i == 4'b0011 ? 7'b0110000 : // 3
    i == 4'b0100 ? 7'b0011001 : // 4
    i == 4'b0101 ? 7'b0010010 : // 5
    i == 4'b0110 ? 7'b0000010 : // 6
    i == 4'b0111 ? 7'b1111000 : // 7
    i == 4'b1000 ? 7'b0000000 : // 8
    i == 4'b1001 ? 7'b0010000 : // 9
    i == 4'b1010 ? 7'b0001000 : // A
    i == 4'b1011 ? 7'b0000011 : // B
    i == 4'b1100 ? 7'b1000110 : // C
    i == 4'b1101 ? 7'b0100001 : // D
    i == 4'b1110 ? 7'b0000110 : // E
                   7'b0001110); // F

endmodule
