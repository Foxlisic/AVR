
// Заполнение данными регистров
// ---------------------------------------------------------------------

initial begin

    // Выводы
    we = 0; o_data = 0; pc = 0;

    // Регистры 0-15
    r[0] = 8'h00; r[4] = 8'h00; r[8]  = 8'h00; r[12] = 8'h01;
    r[1] = 8'h00; r[5] = 8'h00; r[9]  = 8'h00; r[13] = 8'h00;
    r[2] = 8'h00; r[6] = 8'h00; r[10] = 8'h00; r[14] = 8'h00;
    r[3] = 8'h00; r[7] = 8'h00; r[11] = 8'h00; r[15] = 8'h00;

    // Регистры 16-31
    r[16] = 8'h00; r[17] = 8'h00; r[18] = 8'h00; r[19] = 8'h00;
    r[20] = 8'h00; r[21] = 8'h00; r[22] = 8'h00; r[23] = 8'h00;
    r[24] = 8'h00; r[25] = 8'h00;
    r[26] = 8'hF4; r[27] = 8'h15; // X
    r[28] = 8'h00; r[29] = 8'h00; // Y
    r[30] = 8'h00; r[31] = 8'hFA; // Z

end


// Проксирование памяти
// ---------------------------------------------------------------------

always @* begin

    casex (address)

        // Регистры
        16'b0000_0000_000x_xxxx: din = r[ address[4:0] ];

        // Процессор
        16'h005B: din = rampz;
        16'h005D: din = sp[ 7:0];
        16'h005E: din = sp[15:8];
        16'h005F: din = sreg;

        // Память
        default:  din = i_data;

    endcase

end

// Текущее состояние процессора
// ---------------------------------------------------------------------
reg [ 7:0]  din;
reg [ 7:0]  rampz   = 0;            // Верхняя память для E-функции
reg [ 3:0]  st      = 0;            // Машина состояний
reg [ 3:0]  stnext  = 0;            // Следующий код состояния
reg [ 7:0]  r[32];                  // Регистры
reg [15:0]  sp;                     // Стек
reg [ 7:0]  sreg;                   // Флаги
reg [15:0]  latch   = 0;            // Защелка опкода

// Управление
// ---------------------------------------------------------------------
reg         pcstop;                 // =1 Не инкрементировать PC
reg         pcload;                 // =1 Загрузка из pcnext
reg [15:0]  pcdata;                 // Что загружать в PC
reg         reg_w;                  // =1 Запись АЛУ в регистр reg_id
reg         sreg_w;                 // =1 Запись из АЛУ в регистр флагов
reg [ 4:0]  reg_id;                 // Номер регистра
reg         wren;                   // Запись в память
reg [ 7:0]  wdata;
reg [15:0]  addr_w;                 // Указатель на адрес при записи
reg [15:0]  cursor;                 // Текущий курсор

// 16 битные регистры
reg         reg_ww  = 0;            // Писать в X,Y,Z
reg         reg_ws  = 0;            // =1 Источник АЛУ; =0 Источник регистр `wb2`
reg         reg_wm  = 0;            // Запись в 1:0
reg [ 1:0]  reg_idw = 0;            // Номер 16-битного регистра
reg [15:0]  wb2     = 0;            // Данные для записи в X,Y,Z

// Провода
// ---------------------------------------------------------------------
wire [15:0] opcode = st ? latch : ir;
wire [15:0] X   = {r[27], r[26]};
wire [15:0] Y   = {r[29], r[28]};
wire [15:0] Z   = {r[31], r[30]};
wire [15:0] Xm  = X - 1;
wire [15:0] Xp  = X + 1;
wire [15:0] Ym  = Y - 1;
wire [15:0] Yp  = Y + 1;
wire [15:0] Zm  = Z - 1;
wire [15:0] Zp  = Z + 1;
wire [ 5:0] q   = {opcode[13], opcode[11:10], opcode[2:0]};
wire [ 4:0] rd  =  opcode[8:4];
wire [ 4:0] rr  = {opcode[9], opcode[3:0]};
wire [ 4:0] rdi = {1'b1, opcode[7:4]};
wire [ 4:0] rri = {1'b1, opcode[3:0]};
wire [ 7:0] K   = {opcode[11:8], opcode[3:0]};

// Управление счетчиком
reg         skip_instr = 0;
wire [15:0] pcnext  = pc + 1;
wire [15:0] pcnext2 = pc + 2;
wire        is_call = {opcode[14], opcode[3:1]} == 4'b0111;
